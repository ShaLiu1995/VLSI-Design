.subckt INVX4 IN OUT VDD VSS
MP OUT IN VDD VDD PMOS W=1.64u L=0.065u
MN OUT IN VSS VSS NMOS W=1.16u L=0.065u
.ends
