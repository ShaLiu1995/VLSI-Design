.subckt INVX8 IN OUT VDD VSS
MP OUT IN VDD VDD PMOS W=3.28u L=0.065u
MN OUT IN VSS VSS NMOS W=2.32u L=0.065u
.ends
