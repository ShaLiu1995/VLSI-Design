.subckt INVX32 IN OUT VDD VSS
MP OUT IN VDD VDD PMOS W=13.12u L=0.065u
MN OUT IN VSS VSS NMOS W=9.28u L=0.065u
.ends
