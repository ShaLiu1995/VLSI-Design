.subckt INVX16 IN OUT VDD VSS
MP OUT IN VDD VDD PMOS W=6.56u L=0.065u
MN OUT IN VSS VSS NMOS W=4.64u L=0.065u
.ends
